library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;        -- for addition & counting
use ieee.numeric_std.all;               -- for type conversions
use ieee.math_real.all;                 -- for the ceiling and log constant calculation functions

entity controller is
    port (
        clock : std_logic;
    );
end controller;

architecture controller_arc of controller is
begin

end controller_arc;