library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity mac_tb is
end mac_tb;

architecture mac_tb_arc of mac_tb is

    signal clk: std_logic := '0';
    signal first : std_logic;
    signal din1 : unsigned(7 downto 0);
    signal din2 : unsigned(7 downto 0);
    signal dout : unsigned(7 downto 0);

    type unsigned_arr is array(63 downto 0) of unsigned(7 downto 0);

    signal din1_arr: unsigned_arr := (
        0 => to_unsigned(1,8),
        1 => to_unsigned(13,8),
        2 => to_unsigned(14,8),
        3 => to_unsigned(1,8),
        4 => to_unsigned(1,8),
        5 => to_unsigned(1,8),
        6 => to_unsigned(5,8),
        7 => to_unsigned(9,8),
        8 => to_unsigned(9,8),
        9 => to_unsigned(1,8),
        10 => to_unsigned(11,8),
        11 => to_unsigned(1,8),
        12 => to_unsigned(5,8),
        13 => to_unsigned(8,8),
        14 => to_unsigned(5,8),
        15 => to_unsigned(14,8),
        16 => to_unsigned(2,8),
        17 => to_unsigned(10,8),
        18 => to_unsigned(3,8),
        19 => to_unsigned(5,8),
        20 => to_unsigned(1,8),
        21 => to_unsigned(2,8),
        22 => to_unsigned(13,8),
        23 => to_unsigned(3,8),
        24 => to_unsigned(10,8),
        25 => to_unsigned(4,8),
        26 => to_unsigned(13,8),
        27 => to_unsigned(9,8),
        28 => to_unsigned(11,8),
        29 => to_unsigned(6,8),
        30 => to_unsigned(10,8),
        31 => to_unsigned(12,8),
        32 => to_unsigned(8,8),
        33 => to_unsigned(9,8),
        34 => to_unsigned(1,8),
        35 => to_unsigned(14,8),
        36 => to_unsigned(2,8),
        37 => to_unsigned(14,8),
        38 => to_unsigned(3,8),
        39 => to_unsigned(8,8),
        40 => to_unsigned(12,8),
        41 => to_unsigned(0,8),
        42 => to_unsigned(8,8),
        43 => to_unsigned(0,8),
        44 => to_unsigned(11,8),
        45 => to_unsigned(8,8),
        46 => to_unsigned(5,8),
        47 => to_unsigned(8,8),
        48 => to_unsigned(3,8),
        49 => to_unsigned(4,8),
        50 => to_unsigned(7,8),
        51 => to_unsigned(6,8),
        52 => to_unsigned(4,8),
        53 => to_unsigned(5,8),
        54 => to_unsigned(7,8),
        55 => to_unsigned(4,8),
        56 => to_unsigned(13,8),
        57 => to_unsigned(6,8),
        58 => to_unsigned(1,8),
        59 => to_unsigned(3,8),
        60 => to_unsigned(14,8),
        61 => to_unsigned(3,8),
        62 => to_unsigned(1,8),
        63 => to_unsigned(8,8)
    );

    signal din2_arr: unsigned_arr := (
        0 => to_unsigned(8,8),
        1 => to_unsigned(13,8),
        2 => to_unsigned(6,8),
        3 => to_unsigned(4,8),
        4 => to_unsigned(5,8),
        5 => to_unsigned(8,8),
        6 => to_unsigned(12,8),
        7 => to_unsigned(5,8),
        8 => to_unsigned(5,8),
        9 => to_unsigned(10,8),
        10 => to_unsigned(5,8),
        11 => to_unsigned(8,8),
        12 => to_unsigned(10,8),
        13 => to_unsigned(13,8),
        14 => to_unsigned(4,8),
        15 => to_unsigned(12,8),
        16 => to_unsigned(7,8),
        17 => to_unsigned(2,8),
        18 => to_unsigned(1,8),
        19 => to_unsigned(6,8),
        20 => to_unsigned(1,8),
        21 => to_unsigned(2,8),
        22 => to_unsigned(0,8),
        23 => to_unsigned(12,8),
        24 => to_unsigned(7,8),
        25 => to_unsigned(6,8),
        26 => to_unsigned(9,8),
        27 => to_unsigned(8,8),
        28 => to_unsigned(7,8),
        29 => to_unsigned(0,8),
        30 => to_unsigned(7,8),
        31 => to_unsigned(11,8),
        32 => to_unsigned(6,8),
        33 => to_unsigned(2,8),
        34 => to_unsigned(6,8),
        35 => to_unsigned(4,8),
        36 => to_unsigned(13,8),
        37 => to_unsigned(2,8),
        38 => to_unsigned(7,8),
        39 => to_unsigned(2,8),
        40 => to_unsigned(1,8),
        41 => to_unsigned(8,8),
        42 => to_unsigned(1,8),
        43 => to_unsigned(5,8),
        44 => to_unsigned(14,8),
        45 => to_unsigned(9,8),
        46 => to_unsigned(3,8),
        47 => to_unsigned(13,8),
        48 => to_unsigned(9,8),
        49 => to_unsigned(0,8),
        50 => to_unsigned(6,8),
        51 => to_unsigned(9,8),
        52 => to_unsigned(4,8),
        53 => to_unsigned(0,8),
        54 => to_unsigned(13,8),
        55 => to_unsigned(0,8),
        56 => to_unsigned(7,8),
        57 => to_unsigned(5,8),
        58 => to_unsigned(0,8),
        59 => to_unsigned(12,8),
        60 => to_unsigned(1,8),
        61 => to_unsigned(3,8),
        62 => to_unsigned(8,8),
        63 => to_unsigned(0,8)
    );

    signal dout_arr: unsigned_arr := (
        0 => to_unsigned(8,8),
        1 => to_unsigned(177,8),
        2 => to_unsigned(84,8),
        3 => to_unsigned(88,8),
        4 => to_unsigned(93,8),
        5 => to_unsigned(101,8),
        6 => to_unsigned(161,8),
        7 => to_unsigned(206,8),
        8 => to_unsigned(251,8),
        9 => to_unsigned(5,8),
        10 => to_unsigned(60,8),
        11 => to_unsigned(68,8),
        12 => to_unsigned(118,8),
        13 => to_unsigned(222,8),
        14 => to_unsigned(242,8),
        15 => to_unsigned(154,8),
        16 => to_unsigned(168,8),
        17 => to_unsigned(188,8),
        18 => to_unsigned(191,8),
        19 => to_unsigned(221,8),
        20 => to_unsigned(222,8),
        21 => to_unsigned(226,8),
        22 => to_unsigned(226,8),
        23 => to_unsigned(6,8),
        24 => to_unsigned(76,8),
        25 => to_unsigned(100,8),
        26 => to_unsigned(217,8),
        27 => to_unsigned(33,8),
        28 => to_unsigned(110,8),
        29 => to_unsigned(110,8),
        30 => to_unsigned(180,8),
        31 => to_unsigned(56,8),
        32 => to_unsigned(104,8),
        33 => to_unsigned(18,8),
        34 => to_unsigned(24,8),
        35 => to_unsigned(80,8),
        36 => to_unsigned(106,8),
        37 => to_unsigned(134,8),
        38 => to_unsigned(155,8),
        39 => to_unsigned(171,8),
        40 => to_unsigned(183,8),
        41 => to_unsigned(183,8),
        42 => to_unsigned(191,8),
        43 => to_unsigned(191,8),
        44 => to_unsigned(89,8),
        45 => to_unsigned(161,8),
        46 => to_unsigned(176,8),
        47 => to_unsigned(24,8),
        48 => to_unsigned(51,8),
        49 => to_unsigned(0,8),
        50 => to_unsigned(42,8),
        51 => to_unsigned(96,8),
        52 => to_unsigned(112,8),
        53 => to_unsigned(112,8),
        54 => to_unsigned(203,8),
        55 => to_unsigned(203,8),
        56 => to_unsigned(38,8),
        57 => to_unsigned(68,8),
        58 => to_unsigned(68,8),
        59 => to_unsigned(104,8),
        60 => to_unsigned(118,8),
        61 => to_unsigned(127,8),
        62 => to_unsigned(135,8),
        63 => to_unsigned(135,8)
    );

    signal rst_arr: std_logic_vector(63 downto 0) := (
        0 => '0',
        1 => '0',
        2 => '1',
        3 => '0',
        4 => '0',
        5 => '0',
        6 => '0',
        7 => '0',
        8 => '0',
        9 => '0',
        10 => '0',
        11 => '0',
        12 => '0',
        13 => '0',
        14 => '0',
        15 => '0',
        16 => '0',
        17 => '0',
        18 => '0',
        19 => '0',
        20 => '0',
        21 => '0',
        22 => '0',
        23 => '0',
        24 => '0',
        25 => '0',
        26 => '0',
        27 => '0',
        28 => '0',
        29 => '0',
        30 => '0',
        31 => '0',
        32 => '0',
        33 => '1',
        34 => '0',
        35 => '0',
        36 => '0',
        37 => '0',
        38 => '0',
        39 => '0',
        40 => '0',
        41 => '0',
        42 => '0',
        43 => '0',
        44 => '0',
        45 => '0',
        46 => '0',
        47 => '0',
        48 => '0',
        49 => '1',
        50 => '1',
        51 => '0',
        52 => '0',
        53 => '0',
        54 => '0',
        55 => '0',
        56 => '0',
        57 => '0',
        58 => '0',
        59 => '0',
        60 => '0',
        61 => '0',
        62 => '0',
        63 => '0'
    );


    signal ctr: unsigned(5 downto 0) := "000000";

begin

    mac: entity work.mac port map (clk, first, din1, din2, dout);

    clk <= not clk after 5 ns;

    ctr <= ctr+1 when rising_edge(clk);

    din1 <= din1_arr(to_integer(ctr));
    din2 <= din2_arr(to_integer(ctr));
    first <= rst_arr(to_integer(ctr));

    check: process(clk)
    begin
        if falling_edge(clk) then
            assert dout = dout_arr(to_integer(ctr));
        end if;
    end process check;

end mac_tb_arc;