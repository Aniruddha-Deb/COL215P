library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity mac_tb is
end mac_tb;

architecture mac_tb_arc of mac_tb is

    signal clk: std_logic := '0';
    signal first : std_logic;
    signal din1 : unsigned(15 downto 0);
    signal din2 : unsigned(15 downto 0);
    signal dout : unsigned(15 downto 0);

    type unsigned_arr is array(63 downto 0) of unsigned(16 downto 0);

    signal din1_arr: unsigned_arr := (
        0 => to_unsigned(1,16),
        1 => to_unsigned(13,16),
        2 => to_unsigned(14,16),
        3 => to_unsigned(1,16),
        4 => to_unsigned(1,16),
        5 => to_unsigned(1,16),
        6 => to_unsigned(5,16),
        7 => to_unsigned(9,16),
        8 => to_unsigned(9,16),
        9 => to_unsigned(1,16),
        10 => to_unsigned(11,16),
        11 => to_unsigned(1,16),
        12 => to_unsigned(5,16),
        13 => to_unsigned(8,16),
        14 => to_unsigned(5,16),
        15 => to_unsigned(14,16),
        16 => to_unsigned(2,16),
        17 => to_unsigned(10,16),
        18 => to_unsigned(3,16),
        19 => to_unsigned(5,16),
        20 => to_unsigned(1,16),
        21 => to_unsigned(2,16),
        22 => to_unsigned(13,16),
        23 => to_unsigned(3,16),
        24 => to_unsigned(10,16),
        25 => to_unsigned(4,16),
        26 => to_unsigned(13,16),
        27 => to_unsigned(9,16),
        28 => to_unsigned(11,16),
        29 => to_unsigned(6,16),
        30 => to_unsigned(10,16),
        31 => to_unsigned(12,16),
        32 => to_unsigned(8,16),
        33 => to_unsigned(9,16),
        34 => to_unsigned(1,16),
        35 => to_unsigned(14,16),
        36 => to_unsigned(2,16),
        37 => to_unsigned(14,16),
        38 => to_unsigned(3,16),
        39 => to_unsigned(8,16),
        40 => to_unsigned(12,16),
        41 => to_unsigned(0,16),
        42 => to_unsigned(8,16),
        43 => to_unsigned(0,16),
        44 => to_unsigned(11,16),
        45 => to_unsigned(8,16),
        46 => to_unsigned(5,16),
        47 => to_unsigned(8,16),
        48 => to_unsigned(3,16),
        49 => to_unsigned(4,16),
        50 => to_unsigned(7,16),
        51 => to_unsigned(6,16),
        52 => to_unsigned(4,16),
        53 => to_unsigned(5,16),
        54 => to_unsigned(7,16),
        55 => to_unsigned(4,16),
        56 => to_unsigned(13,16),
        57 => to_unsigned(6,16),
        58 => to_unsigned(1,16),
        59 => to_unsigned(3,16),
        60 => to_unsigned(14,16),
        61 => to_unsigned(3,16),
        62 => to_unsigned(1,16),
        63 => to_unsigned(8,8)
    );

    signal din2_arr: unsigned_arr := (
        0 => to_unsigned(8,16),
        1 => to_unsigned(13,16),
        2 => to_unsigned(6,16),
        3 => to_unsigned(4,16),
        4 => to_unsigned(5,16),
        5 => to_unsigned(8,16),
        6 => to_unsigned(12,16),
        7 => to_unsigned(5,16),
        8 => to_unsigned(5,16),
        9 => to_unsigned(10,16),
        10 => to_unsigned(5,16),
        11 => to_unsigned(8,16),
        12 => to_unsigned(10,16),
        13 => to_unsigned(13,16),
        14 => to_unsigned(4,16),
        15 => to_unsigned(12,16),
        16 => to_unsigned(7,16),
        17 => to_unsigned(2,16),
        18 => to_unsigned(1,16),
        19 => to_unsigned(6,16),
        20 => to_unsigned(1,16),
        21 => to_unsigned(2,16),
        22 => to_unsigned(0,16),
        23 => to_unsigned(12,16),
        24 => to_unsigned(7,16),
        25 => to_unsigned(6,16),
        26 => to_unsigned(9,16),
        27 => to_unsigned(8,16),
        28 => to_unsigned(7,16),
        29 => to_unsigned(0,16),
        30 => to_unsigned(7,16),
        31 => to_unsigned(11,16),
        32 => to_unsigned(6,16),
        33 => to_unsigned(2,16),
        34 => to_unsigned(6,16),
        35 => to_unsigned(4,16),
        36 => to_unsigned(13,16),
        37 => to_unsigned(2,16),
        38 => to_unsigned(7,16),
        39 => to_unsigned(2,16),
        40 => to_unsigned(1,16),
        41 => to_unsigned(8,16),
        42 => to_unsigned(1,16),
        43 => to_unsigned(5,16),
        44 => to_unsigned(14,16),
        45 => to_unsigned(9,16),
        46 => to_unsigned(3,16),
        47 => to_unsigned(13,16),
        48 => to_unsigned(9,16),
        49 => to_unsigned(0,16),
        50 => to_unsigned(6,16),
        51 => to_unsigned(9,16),
        52 => to_unsigned(4,16),
        53 => to_unsigned(0,16),
        54 => to_unsigned(13,16),
        55 => to_unsigned(0,16),
        56 => to_unsigned(7,16),
        57 => to_unsigned(5,16),
        58 => to_unsigned(0,16),
        59 => to_unsigned(12,16),
        60 => to_unsigned(1,16),
        61 => to_unsigned(3,16),
        62 => to_unsigned(8,16),
        63 => to_unsigned(0,16)
    );

    signal dout_arr: unsigned_arr := (
        0 => to_unsigned(8,16),
        1 => to_unsigned(177,16),
        2 => to_unsigned(84,16),
        3 => to_unsigned(88,16),
        4 => to_unsigned(93,16),
        5 => to_unsigned(101,16),
        6 => to_unsigned(161,16),
        7 => to_unsigned(206,16),
        8 => to_unsigned(251,16),
        9 => to_unsigned(5,16),
        10 => to_unsigned(60,16),
        11 => to_unsigned(68,16),
        12 => to_unsigned(118,16),
        13 => to_unsigned(222,16),
        14 => to_unsigned(242,16),
        15 => to_unsigned(154,16),
        16 => to_unsigned(168,16),
        17 => to_unsigned(188,16),
        18 => to_unsigned(191,16),
        19 => to_unsigned(221,16),
        20 => to_unsigned(222,16),
        21 => to_unsigned(226,16),
        22 => to_unsigned(226,16),
        23 => to_unsigned(6,16),
        24 => to_unsigned(76,16),
        25 => to_unsigned(100,16),
        26 => to_unsigned(217,16),
        27 => to_unsigned(33,16),
        28 => to_unsigned(110,16),
        29 => to_unsigned(110,16),
        30 => to_unsigned(180,16),
        31 => to_unsigned(56,16),
        32 => to_unsigned(104,16),
        33 => to_unsigned(18,16),
        34 => to_unsigned(24,16),
        35 => to_unsigned(80,16),
        36 => to_unsigned(106,16),
        37 => to_unsigned(134,16),
        38 => to_unsigned(155,16),
        39 => to_unsigned(171,16),
        40 => to_unsigned(183,16),
        41 => to_unsigned(183,16),
        42 => to_unsigned(191,16),
        43 => to_unsigned(191,16),
        44 => to_unsigned(89,16),
        45 => to_unsigned(161,16),
        46 => to_unsigned(176,16),
        47 => to_unsigned(24,16),
        48 => to_unsigned(51,16),
        49 => to_unsigned(0,16),
        50 => to_unsigned(42,16),
        51 => to_unsigned(96,16),
        52 => to_unsigned(112,16),
        53 => to_unsigned(112,16),
        54 => to_unsigned(203,16),
        55 => to_unsigned(203,16),
        56 => to_unsigned(38,16),
        57 => to_unsigned(68,16),
        58 => to_unsigned(68,16),
        59 => to_unsigned(104,16),
        60 => to_unsigned(118,16),
        61 => to_unsigned(127,16),
        62 => to_unsigned(135,16),
        63 => to_unsigned(135,16)
    );

    signal rst_arr: std_logic_vector(63 downto 0) := (
        0 => '0',
        1 => '0',
        2 => '1',
        3 => '0',
        4 => '0',
        5 => '0',
        6 => '0',
        7 => '0',
        8 => '0',
        9 => '0',
        10 => '0',
        11 => '0',
        12 => '0',
        13 => '0',
        14 => '0',
        15 => '0',
        16 => '0',
        17 => '0',
        18 => '0',
        19 => '0',
        20 => '0',
        21 => '0',
        22 => '0',
        23 => '0',
        24 => '0',
        25 => '0',
        26 => '0',
        27 => '0',
        28 => '0',
        29 => '0',
        30 => '0',
        31 => '0',
        32 => '0',
        33 => '1',
        34 => '0',
        35 => '0',
        36 => '0',
        37 => '0',
        38 => '0',
        39 => '0',
        40 => '0',
        41 => '0',
        42 => '0',
        43 => '0',
        44 => '0',
        45 => '0',
        46 => '0',
        47 => '0',
        48 => '0',
        49 => '1',
        50 => '1',
        51 => '0',
        52 => '0',
        53 => '0',
        54 => '0',
        55 => '0',
        56 => '0',
        57 => '0',
        58 => '0',
        59 => '0',
        60 => '0',
        61 => '0',
        62 => '0',
        63 => '0'
    );


    signal ctr: unsigned(5 downto 0) := "000000";

begin

    mac: entity work.mac port map (clk, first, din1, din2, dout);

    clk <= not clk after 5 ns;

    ctr <= ctr+1 when rising_edge(clk);

    din1 <= din1_arr(to_integer(ctr));
    din2 <= din2_arr(to_integer(ctr));
    first <= rst_arr(to_integer(ctr));

    check: process(clk)
    begin
        if falling_edge(clk) then
            assert dout = dout_arr(to_integer(ctr));
        end if;
    end process check;

end mac_tb_arc;