library ieee;
use ieee.std_logic_1164.all;

package types is
    
    type state_t is (ZERO, RUNNING, PAUSED);
    
end package types;