library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;        -- for addition & counting
use ieee.numeric_std.all;               -- for type conversions
use ieee.math_real.all;                 -- for the ceiling and log constant calculation functions

entity mem_controller is
    port (
        clock : std_logic;
    );
end mem_controller;

architecture mem_controller_arc of mem_controller is
begin

end mem_controller_arc;